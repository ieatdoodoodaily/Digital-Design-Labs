package mux_pkg is
	type mux_inputs is array(natural range<>) of std_logic_vector(7 downto 0);
end mux_pkg;