-- Nicholas Imamshah
-- University of Florida
-- EEL 4712: Digital Design, Stitt: Spring 2016
-- Lab 7: Small 8 Internal Bus

entity int_bus is
	port (
		
	);
end int_bus;

architecture BHV of int_bus is
begin



end BHV;