-- Nicholas Imamshah
-- University of Florida

library ieee;
use ieee.std_logic_1164.all;

entity VGA is
	port (
	
	);
end VGA;

architecture 